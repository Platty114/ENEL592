reg include_reg_a;
reg include_reg_b;
reg include_reg_c;