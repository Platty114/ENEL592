//excluded due to my own lack of knowledge
//(I don't think I could implement a system with the vulnerability)
//will try to find this one in the wild.
