//again not a great example on mitre webstie,
//will try to find an example of this bug elsewhere.
