`define TEST_MACRO